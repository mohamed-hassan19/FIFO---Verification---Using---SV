package shared_pkg;

logic test_finished = 0;
integer correct_count = 0, error_count = 0;

endpackage